module testbench();

reg [7:0] A[2:0][2:0], B[2:0][2:0];
reg clk,rst_n;
wire [7:0] C[2:0][2:0];

initial begin
A[0][0] = 8'b00110000;
A[0][1] = 8'b00110000;
A[0][2] = 8'b00110000;
A[1][0] = 8'b00110000;
A[1][1] = 8'b00110000;
A[1][2] = 8'b00110000;
A[2][0] = 8'b00110000;
A[2][1] = 8'b00110000;
A[2][2] = 8'b00110000;
B[0][0] = 8'b00110000;
B[0][1] = 8'b00110000;
B[0][2] = 8'b00110000;
B[1][0] = 8'b00110000;
B[1][1] = 8'b00110000;
B[1][2] = 8'b00110000;
B[2][0] = 8'b00110000;
B[2][1] = 8'b00110000;
B[2][2] = 8'b00110000;
#1000;
A[0][0] = 8'b00111000;
A[0][1] = 8'b00111000;
A[0][2] = 8'b00111000;
A[1][0] = 8'b00111000;
A[1][1] = 8'b00111000;
A[1][2] = 8'b00111000;
A[2][0] = 8'b00111000;
A[2][1] = 8'b00111000;
A[2][2] = 8'b00111000;
B[0][0] = 8'b00111000;
B[0][1] = 8'b00111000;
B[0][2] = 8'b00111000;
B[1][0] = 8'b00111000;
B[1][1] = 8'b00111000;
B[1][2] = 8'b00111000;
B[2][0] = 8'b00111000;
B[2][1] = 8'b00111000;
B[2][2] = 8'b00111000;
#1100;
A[0][0] = 8'b00000000;
A[0][1] = 8'b00000000;
A[0][2] = 8'b00000000;
A[1][0] = 8'b00111000;
A[1][1] = 8'b00111000;
A[1][2] = 8'b00111000;
A[2][0] = 8'b00111000;
A[2][1] = 8'b00111000;
A[2][2] = 8'b00111000;
B[0][0] = 8'b00111000;
B[0][1] = 8'b00111000;
B[0][2] = 8'b00111000;
B[1][0] = 8'b00111000;
B[1][1] = 8'b00111000;
B[1][2] = 8'b00111000;
B[2][0] = 8'b00111000;
B[2][1] = 8'b00111000;
B[2][2] = 8'b00111000;
#1100
A[0][0] = 8'b01110000;
A[0][1] = 8'b00000000;
A[0][2] = 8'b00000000;
A[1][0] = 8'b00111000;
A[1][1] = 8'b00111000;
A[1][2] = 8'b00111000;
A[2][0] = 8'b00111000;
A[2][1] = 8'b00111000;
A[2][2] = 8'b00111000;
B[0][0] = 8'b00111000;
B[0][1] = 8'b00111000;
B[0][2] = 8'b00111000;
B[1][0] = 8'b00111000;
B[1][1] = 8'b00111000;
B[1][2] = 8'b00111000;
B[2][0] = 8'b00111000;
B[2][1] = 8'b00111000;
B[2][2] = 8'b00111000;
#1100
A[0][0] = 8'b01000000;
A[0][1] = 8'b01000000;
A[0][2] = 8'b01000000;
A[1][0] = 8'b01000000;
A[1][1] = 8'b01000000;
A[1][2] = 8'b01000000;
A[2][0] = 8'b01000000;
A[2][1] = 8'b01000000;
A[2][2] = 8'b01000000;
B[0][0] = 8'b01010000;
B[0][1] = 8'b01010000;
B[0][2] = 8'b01010000;
B[1][0] = 8'b01010000;
B[1][1] = 8'b01010000;
B[1][2] = 8'b01010000;
B[2][0] = 8'b01010000;
B[2][1] = 8'b01010000;
B[2][2] = 8'b01010000;
#1100
A[0][0] = 8'b00110110;
A[0][1] = 8'b11100100;
A[0][2] = 8'b01010110;
A[1][0] = 8'b00010000;
A[1][1] = 8'b10111010;
A[1][2] = 8'b01010000;
A[2][0] = 8'b00111111;
A[2][1] = 8'b01001000;
A[2][2] = 8'b01000110;
B[0][0] = 8'b10111000;
B[0][1] = 8'b10110111;
B[0][2] = 8'b10110110;
B[1][0] = 8'b00011100;
B[1][1] = 8'b10110100;
B[1][2] = 8'b10110010;
B[2][0] = 8'b01000001;
B[2][1] = 8'b00000000;
B[2][2] = 8'b11001000;

end
initial begin
clk = 0;
forever #50 clk = ~clk;
end

initial begin
rst_n = 1;
forever begin
#1000 rst_n = 0;
#100 rst_n = 1;
end
end

TOP top(A,B,C, clk,rst_n);
endmodule










